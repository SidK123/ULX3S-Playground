typedef enum {
   ADD, 
   SUB, 
   MUL,
   DIV 
} opcode_t;

typedef logic [31:0] data_t; 
